// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:38:00 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Bj/OzAJAl6DVTPh6IO38KYCitPumjtO4UgGFUH5OH8SRfpTTkZ8J9OSKNkE8sIKu
Jjy4iljB4FOtS8EOK1f6umi75IyAStKvDK89m3Nonz5Lvnth5T1ZnWhz8NmIPxBS
KmQ5gcImgaEgsXzlOYBx61LcDGOOKH8qZNgLZH01LWc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5856)
dFh3/TnofrOLvl5Bdy6A8mFCIsVrGhAaLRnLJKs8hcwoKrcdFGStR8akFzcQvLNg
c/mbhFuTUbKy5aUOzuKXZqax+78zi8al89qxWYsQ3N+zvFhN1eCzhVuRLtcxau0M
L0Y6B66yXidYffCPlg0nLm9lFaOau4CFLCBq3efA3rvTSodFde01O8ZyUY68QpzY
5UJ8y3+0rSRaGoXxIuOPyu3OOqDCJ5O3+RihYRDyHuNT+EI3z30cDLQd6e9GRsgQ
aPNbLs/zvq2UyjUhNhVTdYTIhhJ6FqgwBxD79ukDTTekchsyWQrxwDsoiez+pmxE
tv641BByywVyrYM5uWXDvc+MfJdjm6MRDpt/xp00cvtjrsf7DOqTK5cscoEuVIMJ
mEBS+PMvTAo1m1l6cQ/gcVRcJhNBkjxgurDmLV6MFj3rd8lnm3MTJCuPCXRrhiw1
iNKPWx8Sh2/RZDv92kBdVfZvCa9qVWLR18X1qJRYDXP9NQuzngRcQCBhDr3NyT+P
mJf1Cwzf2C3Ab9Z/W8Pn+FA+HVxiqDhVu6VyFtNPh+plYF9gHpF3mBxCbsRrqZUX
XCtqu91WpCwkuAIHIu1krk/jbI6b2DjpvBSDdnGN8/wjjFn3MSMC0F0HJXd/zjk+
mIa0nW460gAcysOp5v1uddqVMcQ+tedzA2k1tf8mgTm+W75KLs80M76pWigVP8WT
Hxt+lk55DWbcQHrSXFcNuaALEOl4eEgWg3vB9dN7yDoCpdLzKPoiXlcExG9HlUaZ
Ku6tlkZoSqxC7bPOb6KqOD8wIXkW68krE7bcI4KKXqfGK+n0QDNNmQURc3qFlObr
0jpan3DP5l5S9RcZ9KgsCdEId1CvbqK7KjBtfIq9P5K778GbnKz3rIS/WaSaKKyO
SBgsQGUlmMHU+jlcA6HEuvGAKaUHO9O/HmbdD0EyB6XrRoJlo3dB8yS1Ucb1UvyU
8nzEL68IkB0N1Hx2uVfARecUgGEiYNX/AVE8CIRfQeAayta+WR2jRKZUrS15cTK4
1uPE20GIdSqlui4KXPmaki5G5/PZl4i0aVdnrV+OxcL0ZOpVCU+gVnUbMPbg/0pb
wZRfNY47PjRxW1rWV+Yg9LHTmgnHqWsHCKQbh5kU4IqUi5NIcF236P0SgeNCWQ53
b5ZMzmETEKtomFrF8txd3cUK+XP1mlN1Px1t44mgyoII1r7CVNk0e9NC7LBQxWi6
YrWZ4ffvYshYESN0hmmEG/lOIarJ8BTm/wF0ti/95JVEet0xu09E5cjo/yoJi/m5
tKE1QmLdBQh9T+oJka4taJH2hCucIq+e6BV8rR8emy9XR+9HDASKWX8oLNdmZ0CG
Lobu6L8J+9+yO+IxWCz+6pZ3l+PVnkilpNWV7iaJKgiyYuXjQjpsmL1uB9Layyo/
IbikXUnmOHYImYetdauk8XzTOoOSeRI+DTvlR8b4qCK21fqCgfaFVKYSMDGJ8FsL
fpR1cBYXqDYotbKdSn3OqPwUow4YDlPwq9QmngC1Ba3LXrNhRZV+HHcGmatpZsat
PsXxrkj6bF/Ab5GaEzG42C3r4Fcgdnf6EJmUD/AdxNPsaB5pjwVXgYyFqir0s4vp
voHuDKNqCy9nDpTsVcYi6yqdycx961Q4EbDRcIhRSsDd/fyrG1JgsLwJvC7hgtFK
JJmbPMUn4fhIhyipS2ynbA1zKmMPwmlYFWmS73T4xa8FJDUmleep0pWJ5HmOYg4r
2MPFZw10kfP57nhw+5ExH99Kw0j6V+tz55rJMOSfXvYwEoIf0WWT/f4AlAHnvY79
9GVzRRvbHpKKa5nZ0Xtfqgwp+8AAn1ghtUiS7L86RtmrPxW14tNJYs5xR07TySD6
/eVLevz3AoirYopgl0UffEMdUqCggAPJtTmrniPc+O3vV554FjtRhvxQwmsr8Krj
Esbndnfvtfjx2vRfDxtfAZkJngOzKDCbJD0Bb84jYUcchUKsk5roYZ8SF358Z68p
FSwOHQY6sTzCEpIRaJYKbrScXH4pHY/kEFX0aOJEZzljH6zzu3u6b4OuV+xd53IY
CPO4egpRHmgkOhpm37b5wC0zaed0ysSIX/pneXnvyq7NVdqdh1sdo1s7H8OBSUWH
E3QFeVxbE6aYG6ed7tKVcmIC8afeuvmGsJBMjD/AWWzmDsDPAXFzUMMcMvB71cr0
x70upDMSiPijY/ttLROJyI7+EA0FToWnZRgof71+M3HmPdsLgpcLPFaK+OpQ5mcw
+4NOAooAklHkha9b5G1Z5hkd0fEumtazOpLeVYRxGTGEJKLKQTYWf6t2Y3CAlwoY
PxVLCNPa0Ki0OK77sjKEe5VEPGNFSOrgZ9tzdmvLbz7TPiMYEPWy/ZYT9SonfFF/
4uraqn9yBlDSkekSoOiUT5S5mjkoLsdMBSP210UqxLEUMImlTCVJjiAG6DilwoLy
rp7jd5scBr+cc5+jF7skkQO/vKFQgtlkhHtDPizaRqD/bgefZjwPvrNXgw23ZP6k
qArt8II3CaYRgNDWaMZaZVdHDBc0UIYZO1Cahyoxge9SZVYV5HTnyJJcVRzLDp1h
r3wdj7pFogbRe/vHLIJZxFg/g70RSQeqmN0pyEMExDTsH5X+jE/nHoOrjprsM9xg
rErT4+A4kjFfKi8cQyfebrULFHMJSIH5oG48prOi7M4yu7tYnAX60KrGdBvdZ1NC
dDiEx2bMlemKBYtd7TrzpIYylkg5coqVO3/XZmvGfrZ2mRSVz4leK1/q2sG6IE3f
4bVQMSmOemMA+hasEVLKTN+qIznrzqcXMkdO4RpXsWdQ4gK22oPjLDOyk1wq467Z
xdTOGc9pLGgd/xO5Bb0m5ITpmYB1FB9n/X++x8LoH+vHqlvpHveIt3uQ2qM8/Xc+
AjU62yOweNJhUGZmFVUjm4pW84vDroLp3nnNoiybkjwcnc0qwcBDhmW4tLe0Fdwi
7xVwfaWz3FBvWwl+Dfho1kMXpLgwzFUvdXT6sFBGBG5I8pdreguUET+FYARjqfqD
RkpgMJkeMUl8oOwVJIXyedix+uNb1LVULo6agb0844i0T+DNwDFmswTZqplCNv5z
R+DujgsFpFgOgX7a69heidPfYBMMg99HCXQ/LQN2BdDJDegN+rPWJFFliUVfhyKv
8kJ5N8i+T+gAF38nHQ3BbQSbFj7MUDiE2vDXQhBaCdpzAuxUkyipsWl3UEtyKP3x
9pdGWSVwrC6X6ru60zqf0UXnqh1GnQCSlbQC50d1NJSXE4FSqBm/V2DImR1JRqgo
5XvLn9vHsu3xqRYTHPleQoL4eXJmp0DhJcZ8D1mvSJmauuVVSoPIaeYfBfrHO7Dh
ddzq0gwjFhJjH0gv45D1bn/m68V5JQt6m0yh1qN9lAx1KfXa4pwNUBiucv8aRXaK
JPUU1bYMQZeOAg5c5kYGxLv0ctvj8uHiAHjyaE/mxcivceh7ItlIaIHSSvZP/fgn
CHx/NafvREvUFkdzW24kMBp5lPWvXcM1uTnLiuwB0VXAF6gfwXlId9xIW5WoqvW3
+O8YLEJqd0jEKjouwJ2Gnj0AWkr+urDOADITAGZPk8rAJJwIDIsfJpmZZ+EjMHUs
gwMlxbxMc5JpCaPBDNqG9rgLYLAvsecXWD+FRccpyVFvJIRv6o0xgwx5DAJ1m8Ro
mAVdAQ0VyCN22ueju3n5iBIGD1+KfzzHQuWh3AdSnXrOp2DwlADBG9F7ksoog/VG
NDcQw/NHky4HvVFaSz8Pm8wKI/uf7a043BG40LkrlO/Bfm/G5JSBkqKeH9IR/CUB
NosdTMKnVqVvWGkuNhyVRI5ACYzlKbm8b7p+OWDeSIcq6l8vLBZOF3Rba0ZZ4baX
N2RAOUT3boITStHTbusk+HkBR7hJ0Pgsq5BS8kk844YtgBOJM6WFHbRBnJHFpf0L
c0tM6iLSZvXCiCTN2i1TAu8u9cx3Eo7jvv6I7jrUbsVeOHZUMkBswJwUBN6nsL4y
QyiaRf/GQD/rbDXxCV1usj5I5d9WqDQ0kIpOIj6wioCAZgtIQZ+QVcsX+nzXuoLZ
xxJI7QF3BuGWGDG3t+e3X2Ty12OE3o/VJVEKXeBS7xlDfZfMOf8I6nYm+4nev7GT
upLealrMAmeuOCGMnx33Vpb1lkGKq33488BPdgTV94gFBAA0VtgReyDHUXk6VWna
D1X6dfdmJeWWDrVV8jqd0VTicebzzMyOxKYf9FNBD9/TuiGvlf6cyn7oDXO7ZldF
Q6BybDkFQgq8TUyoMgQjuxx/OmuUEi16ZJePnI4p2v6jJHquHvp6HUkKVOvg3BPO
xtO2ure9SEFaPfeKqy+gfkqRILIibDcBz9BuoyKMqKceJ2TLcx95hVR/IJxeHTP6
n6zByE99StkO6VrAkxc0pgpoqcKcbMfcIHelrb65ORAcpj1ZpzzimNfHnGo0UFG0
70TS+46ebz/Io0YsxWC9yoFJwA2EoDuoJ+CdfnjCH+VUmRjSsXArMFaPfXchdG9K
xTPnDmgXGqsdtuf9B8Lk0JM95efvx0LFKj8MLkRIDrEO1079yjmnhiCjbw39H8Su
++oZ6rKlV00r8b4D3twJFEmQ0DFiflXyCvPvU4m7fVNP1SfAKkZUXV0VdB/swC2b
LQVRWE2ufnjX1WOiCe1eAKWf08YLmeLd6QjtHpIecLEHazDZ7mm89A9XjcHnhMKp
jzsBknirpAECKLxGvUi+apmSpqJAHW02UnkcgcD6NtS1tLLn1ySrWAo1/5gSW1PV
5GLMpzua+p3o7LOae798m6IkMb1SVsjrYBtu2tvvy/r+ZZTdREJ2pODzOzeqkiAq
K8YVh8cVG3ZFL+IpT45W6YC8SjYPU19WcTIrPInBAKJUL6IqTlX9b7FmDOYNXtSZ
1ViALt1AObstZreFclPoO5785KArXzk6s4w4eVU523mqgjtlfNGmL+1scOrH62ij
aydlrBQQOvad9mJ5whFtB8AmX2Hte/GIqoaPzgYpTtDrQaQBV64HK4GX6TwcFWnz
Si08eHGoN5VZ1huqkjRffjov5iudR37dSMyJPbEvcY58YyV+L/N/HHvP5lBg6xXz
4z1dlNk/YvLmIeqo0jDOgjGvcMeELq1+FzfiqX0ikxBugB3fXFVuSQiqWthpbLOe
ojDl7R0WRoC+QVqkA9ZnvDSOKOD/GslsFPb9Nmd8PMAnWJodcyiBkc5wpNe+9cQv
508sLTrn+2GuiqGP+SuE7s8Fs+b119nAhbDAz+BAQn0Lyem8IohFTO3LsP2faH+M
vDZBQu7wRDDEuzBTQyuL9BeT+DiDOD27bNdBQMJ9Y98v3QTHZUR8IARL7qfNdrQV
/0dgcG8Wz5zb6qN8DDYLWVUYxhE8AAJ8BtBmeNeT8pcGFQ0tPFXa3eAMELu8Ys9Z
C0B3AqMPVRJj/4TSTbInM7eoosVUm4uVohkHvaa8NjyHbbNFjlz3MNhsfWAhvQ5P
f+8G+WVkhdg+X7skODa9hy7hwldZxlBJqbn09p5jQKMPcvXs246BBtYNXicdlc24
6lt4x8p/1KdI23fmtM1pdCEwfTtBBbdTKQsNSkvPXYbuj5v9kKGuUVwcl1HTvTA2
gZU1FMGcJNS2xPjS6E3Y2jig69mVxkYDxcvgbfgtTIZMjaDW19E65uRw1k+ktRW+
MmOuXDSXM7I0mpzmM/fVcDJbMDJL1x9Jhfc7o4QjPLnTCek0n5IcPCrmvdnQittk
DaHrQGV/9CH2unGmuOTFEtbt/OKjR0txuBfVsrqyXbIQoWsLIoVJKA0N9ml5Pkyu
iBWdbBpqcW9ILEfJVZXIUlojbjO+ym+IrqPFzcMh6ky8gqWbVHuFAlQrQkTvynrN
FRlZSidIkZ05/XwDkBCYhwdflWG/j1bZ1yDyU3aNZliyiymHukHImjPLkZrw5Mo0
r/h2A4Vp2OZYYzxjiIgFxRu+5VCSuIo3eRahB4u9MOwIRuk4DSKkw8blQoC8zbEm
hGslFRfLfwKwAwDytTHDJhZuEimWjtsEBo4DA6dzPYPhhYkaEfsxQqVNXpYqqLza
IxqgnXZaiWbNNiW4+SVTnM0Naym7wE9i7fMLvq96SWewVvUlqJOp6EPCXMw+6GEu
JnO8LxbJWGcxyZkl8cE31fr61gF4x3GaqqS/1NPkhscP8++SNtZ+9jaVnLK6dyGH
mUDG56B+vJbw8up2AgILs6mfNLlJ79C3dA9QqGka0GcwcsIGHd8UGr6/Ba6bgkDL
xOcazqrCuEUCZzhs+rv28hHjS/HH+1seWF3X159EEjdO6NPNk1JzvOE9NcfVg0bs
4dhvs/tPetFxPQTbSSvlAfkgx4PQVXeEv+TpY9AkqEYW2eAQu/kGUybIktefbpEg
QXQAx2lthbyKae6dy0a97nZmyKp//utpCcgFzZKdgNo3wbvp3q7ZLsU/4A3z34vU
M7DDuquvs3AQeZ3pepmXebrT8xtuY+dj2WiwHNjCVXHFfqKtHsnX4Wu/PEdpcq/3
2No2D4GyNAexNCR6DN7H4J+ZrC3ZxvbQcIYvIf8lbtKVEQeGks7jDxQRC7w4C5EV
77QzDLAR88VsmjAxnlBpeAWZD04b3HsTKxhdhiQSEy/TOwGKQjbTc28FGLRWjqSs
xAeU7qDn54BwKC6z7XZkTJv0fpomEnnf2G0oGzQBRpy7zxQaH29bemEYkal7VgIZ
QDIUOCgg4FiNUz+VZMPpKp0WSJ2/ZX+HuYTVgia/PLulnEhNqJIboMmpHBSn6whA
+JuLuomnUYABG99KDdRZi4GaMtxtBNBUj1gcpAAWkUYrdOEIHardDi4lrJTfBMfu
ERdFG7KakDopUjQWj9JG2j4HRitVr922j426aHq7NcJAjU65s3wdO3p8T/QcwoeZ
ob+Uh3EpKWRxp0rAmFSESrumZWEIxyldIwYf6ctyFmZbQlzrE+w5wy2vsxedLjlx
6G6yaFa95tS7xcx4zLt/jd7r3ncQy++YrqomJzi2dQChdn12RjEkFohrGxDNZ2YK
lFta8HhXLowR2aoUbg1xam48Lt9wl8+nnKJreODcekmD7toVxRenZF7NvKBNsjfD
FtxJZaqNdFnrLsQmslYa4xuGoAvztt1Emfy9PPnyskVzVm7FUUP0YkzfcKuumcDa
6AF+dwGgLwNDB5yyPH3PRXhYMFx/inkagoGtwJpFrVhps6fpBOwx6VLdCogU+jSO
9hlQbKcxDxciZnJYQUYpdM0fmb65/GNnxVLP23f0Pxu1nGWopKGf1KrRknCCGTm6
Eocm4kA/b8jMJfuZN0CmqQGV5uL6BqicBlo3pK8D+KJ4N9tBFJ/17voBU7VUHZIh
nAKe/RdmImgGeJHqie3XUuxxfWUwTwKTwOegQO1WQCWIdN38uRdfBUvWiM1Kgt2n
XtuTFrs0ZHTJBb1EApzfODKC+VKINkaK03LQxz4Lrt0Spn/TSTr/sMkMVpztxz1y
HGhmVbYsW+kJ4UVJzYRiCNucrH6ROTmt3GeZ4mHx87l8IwdbLdmqfRCdXX0/WEGV
FDTSn+k9Rp5pcU0AY3dscG93ZZlmT2pWUAYV6nLOVLK0aK8VAcvrjIa6QyiUVM/0
HaXUY9AzrsOxdpO6t5OkHR06ttsxwJE5bxwJMEWe7OlGfCcIpkhyOnwjgtVUPrBC
/PUq727wPMV5jlO4fx7f1RIY8Rwjd104/NT7p9+f53uUkPjsiWt0pBBAzANm+3Wy
VqDPcj8VrefA3NtMmWOviq711IBrTDWB9x1Q563SyMskZOJLulwIVt52AfjsJrS4
M/3DpL9aaQJJXO4Ju97roipFI7VB61TeUSZwmH7pMFU7wJbFDgZLbZpzndZfOSB/
`pragma protect end_protected
