// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
NR2PienxwY6UZnzOjiUA3G68eNzjftYEQN9Q4B4ZEa18Vx6mBkMAzfqwSQ/8eMeune4D8Zpp1aUH
ush8t5xgADuYh/AiEY0CPxwzx7cC8VkPZbPIpzCDfoSa4qS8DGV97ZQiV5b4V/kUJArOvXrZNAvK
4DFE78odSNpICvmoVN+wc5UXzLe1UuP3MXuZEFDFCGD8RBRTfwfkzfKH+YhIucoRjq33p8F4WoDZ
99aK9TPkWpZ3aiGOJpIFz+SfMXMza5sydTGc9jlFmeyl98AzLuSUw7cc3uIDZM6Er5lGhyAX1jvh
M64ipRyHAlc9rnRQFUVm+d3YF7v3o9TvydafTw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5264)
IKnOyjX8g2oCRetIM9mNVyn5hZouFHyGowEN4t2XK3ySfjyhSgMypn0nUdoBYE6tV5MtdtZlfvDK
48W+Vlj5ZR87iKYhvZMRGILw9FjLeKq8CTuC7wThojVSV7GstsQEWya6weMbOfUs9kyjKK4rOeOq
ryHEA84xJRw5AsqP/aOKBiaDvGI3yXNIoFceLSlMrf0STkD3l77dW6W8vyp8gjk1NOAAh9LSADRu
b0d7HKHiIqWR1G1CPLKxUvCFTNhP9OTD1d0TQa+0yd0gYJriquNUzyW6rwOIo35DcHYX0NDRi4mw
LAfap0MEbdvl2g1cS24RU1oWDi4yw9QMfGBsbeL0P2Gh6cKIHp3xLzEASbRxxrlFXAwkEiNmPbHy
tq14z8XexPjPxKXjaHteyNRT9GnZETyP+o9Cj+4x8Mi6AWSJJiPcjGoMCKepd9eMG/HnOG+b8bdj
9g3VwGIWcgTl+BcVQmlqs39V87im1jeBmOP18IvwzbjT6FszLXMqphRD9S5DaAhy77DdrK85Djor
z14VIZe6tanU4bC52rRNhUbSSWM37xKiHN4wdtNTNE5/N7jD4AEb/zZcSPrFvwqFY4Sf51KGk6ll
dLvU4liAAt1cUx/LbQeZxjraaKOLSl+tMqNwSMHHBwUEjinoQDi36Ubw90qzyLcMjPgfCIwdbWq0
M4FzqHJCRLmSHFWddTJGiaS1GdeeE1koJtjgRHVP7GPhCdURWW5OYftnJPw5u9xpM9UgNpenYNQ2
mmyE9L9mo3QJJsHnfcO1AOPEsJktnO+b54v+w/ppYHSS4n3uYjH1tSiAK0C/Pv2S7ppx71qDQPaA
PaNOeGwqtFTgpDVMdpOugHSp1Uj7DBSPZM0uN+ervOl3CIX6tCmBmCT/Vchm+iLXe3fekltk5JN9
gK7NfD6tvuhAcyFCVqMjmg8cdrFTtZnxMvMA1/jstTkuCWf8yZs/i+VRtQ9+J8Y2w4TE652qhkoh
ofwRrY/0pNXZaGj8wRdHeXWRGceYeXaaiUaV2RDcS6lSpJkkT1+Kdlds0cER050h606VamxYmvgz
e/sGQZeooyjlrZHzIjTPyq92q9fV5GZ5cg06gqyyXhHdXHiyNbh/wTkq7/B4jPWK3c/Vfyg/DM44
KnjmXotBa1SZqvyw6eR1ITJaFXh2Z1FsJhvxdk571ADxli2+eiXhlpceUeHtdm/lqPOcLrKQboCv
o1w8qFlJJCL9a1betuhhgG1CI/icPeCIH9JPOh6Fv+SiOozk+vdkXBgtRMk1u4v6oOtyC5gYGB55
ZoNPKveCZbqrGLysTC0WiM90EzCdnHYd407No2TtdjhDS2NklpbrdjtGGnz9z52SSMFejA/6Ld9A
BBNNgmmtTlhgYmaM2/xwY3N+f/2/c2SqXziDkEIGPiVcT9rerJik9CLlJcqn0yU9MWEKVYPseG4g
mEJ6iLdjVXTdGnR8o/LLASw0clyQeP+TsxfXeReKCTm3jGeE78QGFXMuHgVWVA+StPbp9BoM7lQp
KsRbyYrYCAxACeUnWUSMqhvO6baBJBOC4djbCMN1D2X+oQ6wM0jtPllqIdSAPM7CySNb9kShBETe
rPVD30WqdboagQI3Wv6lYyszcR0USOoTxpE2anXouR31VXlcA4cY23j9oCcS2p5x3r56rFV54wNt
IvL4uxcbb3Zige3d+9+6iR2ZoOWfy8lNFc9xPXGlFY04/5BPhsUqVRY5djdbjmMVwVNFI6dl1Hmd
pupBdjQ4tSKSfzPWoRTDMN+VfnwWE1CETuHpOS95xEfTDSbVMWQWopdX/4w25++NL33UUHfEid2y
555xD4pjRNUN2xkhVYoaoXri6fNSjghuoK4OXfhwPCvWREm2ISGbmsvh1m4JE2G4EDEil5TFmK2D
DP8RK08bT9soOIsXk1H76/TRGF3aFXMTYPARbNKndOd0TyU+gGKAOKPwEOPuyeFkfRvJoam4xmwq
6X5015XN7XjvhTKmoEVa4PkWUziuV6JpmkLgmBmBcqIlM9eVmkUg9oXvrVnmC8uJ95MWnk5dXjzs
5Skrpg9yUgntTx+k9L5l7WcF1N1zj8HBIpV1d+aoJ8lPst+aBAtVZixLMPPLuy27vMr6gvZupoxb
D2rl8DxHU15OTPE7ehK+/RSqSu49wlqZevswVQBO3mUvPsrFizT8f8Rx9K8tvKei2kIWz4PuJpqX
jB44smj+Z5pfF9yl3cbe0jw9X4maW1FFQdCnHoGyFrVkCcC2plQrOH8wtXFylYA7zYrtDXRbVZrl
XctSRepwoy5UOl5XX8XxAstIEbmhnHcQDsBdlIJXSjDXgiB4ZaNTloo8u2LDK1EBP+NKkpuYc46+
HUzUQvy6USB7S3fHwlsh2P9H5gnr5EDHAKd7zoneRZxX1pMsTygAkhzlhVMlQUi0PxZGoZOZK94X
QWw7c+N3gNOqfKLVNU02oFOMpFuu40CLJabcg9tHqGsxieFMx+o0D1v/h33tfoGH9rnF3Z9PfSJq
7WgWFFosOzU6X9zJ3KQGYVM5brMDKbPXQMOhzJ6+XT8Ie1SFB1e/P5Zev9/HbIH4Du2a9+Onu5Ay
68uZTOVooSIa4DCoEkgllzEtGIyeILCx0tN7jYM3s5oO8h8NnFscvymFK3yRTnuBoqDRTuE8iJIf
PazBPNgJHrmW1dJpfBp707lDeI5xPki0uGSSbpXt0HJ1K5ncLoW8nQlenfXzrdNuC7ET4khAxteB
+usjcdbcL832klOrbEw/PBj5/K0uG0UGRTO7XVlQW2k4nZ5lvYwvS15xx072uE5GdDe5D74m1biW
HGKCLR2EOrQEdVmijLnWZMFaFwbVmASacA7k8VjuCcFk17AsFKxy+9WtbvF3DS7BWSMpGt9k4aU8
rSeC58NF0G3Itu2jCWP/EFnI5DzXfLN0Y4yXUzgM9X4hUYmawAW9IxBGOae1WzTWJJ0dNONaOjBi
65i/zsY1hc8Oc1wfHzJ3HQGxiZ0i5J0ZA2/Ienq3DntUhCSOL20fZjTcwSRz1NPu3vItM/B1CUg7
ibRMg04GwOcEoKe9dcZzbuisRzMtHS6xABrkZZXWV/f4bquaj9/MoL0yXNAaUyqDKWTC2XURMy3t
M+5uVxlH0auhJmC5NhABkFbjzbGeaDNIEFk4Yb70B1QkI2qwd/DcFr+863ZEO02hYvBLS9kzvHWn
76nkQ7dmBDSX5exjBFVtPat/O6HLvBz2T1uKXELamDNlZbXSaCtqWx+pMh+YXwuLSUq+uy0vKpjC
hRm49wiIQGfjFlJwMQgLSOYxutwQTIDrux8VS5OxjvLtbE6YRlTmg2QCHpkRXQ3v4IDI0/T8jwyO
0jvg19zSulYm3fpCfTe8/PwV5PAd+slSpQF/6EP/WaZpAcuqlagk2s8gmcjIXqXnYWXTJO17L40V
DUUdf1zBURjF0d2YRz47AfLf0msbEyTbEdP7ui6TgAz4Yhq+wsMT5a/XxdTxpy6d2MXnph0dpHuq
6YHNluRHIeiJd5RU0opfEgnmrlYNx5slilpfXaDLKdDQTyUOfbHcGc84d/LN6+yR4VJZQ7BUtUKH
9UJ2OUTKefxCh42aUGZxkSWgGsW4CJQ7R3pHJOt3f2q7HgmP9+ReFDwJZg5X+ihNKXAc2YWG2w2x
s92RucFKLWgLWKjvB3uCVgbL0a7EYzWFN3Cm26PSx0pw2CHrNSe3VeyIDoUiyKMd5nlHLA6vjfDL
tGlwLM6AYTnc7tNdZygq4OCU5idYWTmW4eUMaS/YCd6ohj9VcfLyXh/5TdzXtwLGAUt6pUrxqhBZ
f2wpx9FXIyefyQWJKCpaCcoW5w9jeOGCxlA4N6Zjb0D7disdl9f4xMgfH1E1Rh4HzLcMcE5/HwQ3
ruRMdn6WUC1Cp1NubnV5bAZgYQW9KBhaMztKOmLP7Bm5l26gHQ+LfiU6nlrUfz/xfz/aFooTV1Ls
Ngo6G7CPn42QxemC1epCvPXO68/sW46Xw/saecGsIAsT1A98thNsuj3t29c+B07Lnopj4wy/9Mp5
C8P8uy7K+q7CNH5OMbznKtpUr1M7DJP8hYU04+mdFXHh6RTbeEr+4/n/klCKfyVVjvJsAmZ4WiHC
Z+wgmHBJJMPG4HIrmKuVAJHvvdwW9NNUuJFP1wUZazaWXbUZjSYykQ2wkN/xdhYXpJpvhdlNcpre
1AnqtRVR2De5/k57+/6rgDDz5iCG0Qi5zBkA1Ku2Qz4lk/Zd3SQ/19sGAq/o3SIpfO7lvcqpm+Kf
fgX1UnLj8bl889J4d9ala+yjzOp+eCyFv7BNxSiq9cVWXQYFrhcgv19jhbFcwVhfalO0iWuBU+xB
3GGPa/c5Y6JVBF1SgylB1VRgWgRKn+AOqEQvXYVj0uI6N4lzrQYh7Tdidw6oYqiXgGfryxQtd9h/
B1NjgmskX67s4+PDBJmbpaFeeUn26gI9gwh6218GDXgIr5gWyIFj45EUAyMDoCbYn53zEh2zXYaH
Zxi18K9eDj7UgOA41Jnz+975lRZPPC0YChpFN69HtMc5ODyEzkzQlz6hpM8Yq6JDNn+V/uRMPCUJ
IiLHN1VGDWEwqix28SzboHJiTijgGhBB5il++1hS1Jqy5AAuSMjUbBFCW99ULrNDS482nuKJOzcK
pdofrUfOlOXVPlS2B0ODOUO0l/xWQYCxvgJ5/MPBTRkrd9yFpCorKvGoKN/j46J5zNwzP4bx7szv
2B82IdTSLNxAzQYD1MyOcW7BRoWNHNeDP8rC454l7sn06Vqz//i+WSYHpzgUbey0zoX+19CnkrW+
Sx7pRUDyPd3h82fAM+WaTRW8l+x8rUtHpSu2V/C5bSVYQtLPLQH1RJ+M/CJbcitrqxYiqf/xDuOs
Ys6Nv21Vpw2xO+PSt1vRWZCnIMHFELfpxCZh+UEyHgofdL0aImbq1lFLbJCCeGYhW5/65ynN3Zov
cpHjddESRWhiNGsN85Gol0BcQQVtZA8aP9477Qh1opt+bagCEDF83Jsymf/jlb83mivTNx8lMb79
3TXgVODp9bfzKiY9rUqipkF8iM+r4xPCJyilfMnL3lx6MZxoQ2Vw9Ikz1z9pwQYQY+0ETbasFE7G
QloQ1hQntE1TxvK98N4eIu6x2qxZRONq7gZQw5puhyamS9v5OUFDwEkf5HPezi05z1N+cZX4K6qL
nnYK0l4/gtG7IgCz4aliszOuyu2utAkRZn+8g2kORi93nLDX8PRUlYhT50PRDTykyoA4eo5FmUIb
+YV+azYIXs7CwEwOniVQ/aoxrVrGx38cGjwWQF+qabdEw4NZi5FMr7BWFtiFHUic/r9JEmRsYsmk
jXH1O0HqfKSYa4s8HE+pEIn0wiFfdfFR+Q0vuy+7DABfqzgv5rCfXlshpoYIBuJwtv1dv/+9Syrp
x0Bur5OqpZ/CDtaWYoTBpV5m5c4/T41c6OsarhJqi6kpN2FJC8qO8VDgTRON+quiAoMFWsg/1JTc
dailyYWsAHA4rpcs0gHzJK83EykCU3H36UhX+hWo7g/5f49VGQ+NyAfeRKzS7ipUisA9dV+KmOdu
VChhMMh4f5JKWvXo6OFCOZF2qyj9iiw2OT8GbGAP21PK/txPdMQXJU9hz0iEld1URm7K3VkSO4Uy
GY9OaHYNo30PI63QzgE3yJKXBRtQiXEn6UlNmUZaanMSYH933kzONGQGFDh9UY2RF2xZTvxTEuI7
kBQyNajbl7ctGScH+fJTsevcM/IGPe8FKtEfmO2eCHhk5bajoCkoozonPq6apQqiWhYLDBWOI/Xu
s4AoFdFbzB4RgXU6d546CYXfGNpxlrPTvvsv++nwCjBws+u4dwHxh8QP9rU3Vqea5kQSq12f7akx
TD/2HHAjcXukwAV7dRnL+Z6GUIl3+KG/cUq0cLBcg0xpht/I1ldhb8l25FbrsRMD/X0x65J+jy3p
ZADY7km2+W1aIkVzw6PJxKEsBdEtCVOgJ3uzvFQupGopbUmMa+4kj5i0KESSMR7owFmub+by9NFU
rvlw/ILzB+al4ri/24b9kPpXhbFeUhaY6LM8iooHrqedNsohLyc8LMhSPoIpkbR3DtKXuH77IWjx
K8GssYyGD1B/l/UU/nFxGMpeoBq8uP2KvUJ2IfR6+zBFhxlqzqVsORPhcPmHTGzeO/Ah8b7bZXd8
owgELbhKLrrDaZeD7sj17Qz5WWiVww7LUYnM8wH4Kf7luNq5ajc2AbmTLZODjXTxTOSEsGVg8/7E
MhW3BlWZwqocZa3BOOkQdRIclIda5N0lzRSJBW31+211IwyaYrvq6IEYi34JDgskHSM37wReEaOn
9whhq9EHYAbcsEykV1IlWRjX/LYgkM+HhONAsIrghm6y7fRf268sjEbF12S64Kk6+eZWlJbJbNR+
d07TgB3i6y+jnQIoG4/BAv/fpbz93vC7/8GQM9kgG3tKR9tc0w/vrI8n2HnlRCqnF9x0JITkeqlr
pocExi1Fm5Jhta5bm6mBLqpH5ttrccP6ZahnV4ZkELp9GaJmQVaSTbza2LyclS1mXAic+scRtu/5
HxBCmyNs26powScXh7rZLSPopIBGnx7lcEh7se9DdOunTuY7FPHYhvD+vdvwmS3FIfVjOmEwEJRJ
RKL0cHMUe/Z7xwLr3q4FLlUtjsp7YxdPcyDDyRgw3anpoH5oAtXTRpe8oF3YBndh/KdGCPqesIpu
iSxFbbTP3M2Vi8c3JK7haUktHwwxP7WyULyid7/6eZhvQRGmOzCMW7ktN+CH1ij2aoLsIkzYMVAT
JjwSFmBO3VGvgEEc//jeoocTur/3V1hkKFejjKf33B7ZhzghByMaJE8gKH9TXT6RDfHH2jgKJfHq
DQhygkae6wVI0BwWEjD806ahm4GvCuD8DB2jK7p6V0GCrVvI3rV2KptZpsQoHOITJhAwxm7BCgbz
KPkKsNvKqdyI+64Bq9k/kU6qQZx8ww12YdS/apWprcuP6J/NfRURzT3h6TW0UjWB20a+dR9+ATob
VFpj2/sJ2gTWpiI5ER1adLphlUY=
`pragma protect end_protected
