// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0std
// ALTERA_TIMESTAMP:Wed Apr 26 13:38:00 PDT 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XBSGpMZVbIt1FX7K1RDyEkEumec/VVd8OUrPBJrxXQf/fzF9XfbUM8isfccqbcak
l0UPidVdAa1PpG3zbt7+Nk9aoJ2KQeJZ6v0X0peweTc2pWjUyKwKJ2jeiU8hs7CP
Yncb2zQcARUybiGv7HbBCyvOeLIzZwfypQ3y7/I/uS8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5344)
cCELYdrTZov9IneEBQIH4X4mWT3pz/VHOg3URPx2IMzs6XHcOOEktYBWdX6imRbC
Bc26rYu5ln8qqA19MDFW9A75R3yRU/I4z/XS8aI8XkHBXKmXkJiyk+nxyGrtGsvy
1pzzE0I8xGr4RfmoxLlve5ydsrmclhT2hTTHDrV1A4kLnrRW5+VT3cgot1n3Sg87
C7G1RggKG8llNfqHX6BS2Zf+nWnvlaSr6VrS3Jry9WyFBnFAL+jvrh+EIwNpqEkW
d17PKnRtR+G9mS7gI994eHWeEZyGIm9m8CCz91OPuAJIrWlaEL7RAvXPOZs0vhWf
xa9x8XJ/hIyflK90Vh2mZGhoNLm+dL/RJvFff2E+40p9ICNeVjaPRlmrzVOS7J/S
eKpMnDYPl95HdQC91NvS5m6S3v2hTx536R/0kcb8YpVQl+PxGqxjdXjQHkkjQWrS
UCsromQ5l+EZ2j6jmJqx2KadrL/Py2OHCkJ/CK2WhWvv6oXg3vFidjzSO+BfTsWv
hWuDr5xbkCNN3fVcgdT/Wj18Y7X69BqNo1vceLI4fkXJ0Va8mYQBEkwyeauooDLm
2dyOj/FXdIYBCeTr8h91GzX+5YVGJjIe86OtuBs8QwiBG707UCunIU5ASGlLl5Ic
MFAMiOYkdkUh3N/DXKk6yGf+W5jRuCLrt0nv5dpk2Xsx2/j3oCn3RWKU3bLkKEoI
lTU2BE9TpDAHD4TYgN427sk9/uvtuN3e3NmsXPHBgfiBndTKc14s9ZEmF0E2hGf9
US/YWM4FMr/D4NksRV4XV2P21UidQNIKwvhxhFyz15SExR0cRhHspbZBHfxFkopT
C1jQ+cdvRv4T4xC7i37fB6+xG6tULraqDI3wTSSslYVNsBekOrFIp+qY9zLufajY
cg3hbzHsrwUY0YtM2UcZ1dkfj4t27I5RCJIjr91G5ea63YexASV1dWHxX/1McgH7
RvGz99naXd3trGZJz4uhVLRs4k4EbQenk2YI53OEnGrbJv4pESehKi0Aacla1fuH
qlOw0/rt3Mqm4oVTXzSCyK4NhuCyP1S/dyjnZkqj6UvC/t6nE7etnphGBx2Q6ZcD
mGG1NKGEWQJADn2Ju6CMcTxL+03jGkG2colcscxh3NmZQWVcRF6OvcZngX6H2qS2
slb0NJOQp5+Vm5qMyXhLZyDq8XE/XObKLGMcpkH3xZVY55VYdsb0fJmWqf4KWakk
I2ChHpsAY+TDjkBNrUN+VIfAO1W1g+wTw6XrSseQC6GF1yLW1DO0ObTDRprCm2jt
Uy28aIs04DEu73PTtaPWTxJwA8xVHO8Ie9oCVY+ici5EexXQyQ0qao6bjeKVU1dO
ZCL3CMwIIOuhdvtDziblT/HdI1/Eq4cM5vtYOue4gJOw9BxoyCeSELm74JJhMifA
LDeOfK86H0lyzP2MqeagiUiPVgK5PMpcNKIbzpLTPtMtA78djJVy0xC/NH0PGX8f
al2v4u+/3zyJGLQrR2bUxvGfOmIhS4HKz5JfBdNMLk18b3d04EPyigZAobv2KjpD
iCp7dyVXN5tNQB8sB2mUcukmVVP0j2XWd/LwhR7fxgRy/b3lDMi18m8yEGr62Wgg
4wODWvsRdmYWhUx4aala4GAahKULmzUG+Das+cnfEemE3v09P+gPm521eCECExY+
4Zh817nEGdSvZRnX92thZqX9fuSmWPgw4FfbGiWRhxZHEE81zoETmvxfUj+3Fql6
YcykEb0Tu6B6WsBKt7yHuSEdLhDVVgVQ664Px93XdOmL00IVlZxMKh5llaNcTOeS
rqK7+62DqYDsPbf80Jfs1+2Bp3QGFxU/ryYVJN0yXMh3uBtE4ethnCHSFyFtBotm
hIqcYi4YGVg2fELPCFZVUyoH88B/mHEpN2Alj6JVjZHeIlRc64068NjIrQJAxHhh
0CVrKSwxhsevoOvGpoxzSaAHACjmikdWQEAuQpnB6BZUXkNjl6kar1BGqyCvKCmd
IDRyyoVRgtzIfMg90tmz7atp8/Gu1HHNVtRkNvPST5K19uyITrHlT4Xrn7Mt6OyN
6/R7SGNXGmsmF5XfEztQUVGPRk7jRoMN8tiNYlN+RjeHshNnisid+BkcsHuZGRLE
z4fsC/GRaQfd4Oo6cRPAKzy4Tcx9XRm0GDX76FkGYAvRSk2GAjW4JWHXk34j8ysP
M60JoJF4D5cFNMypDb3/8RWcR0hmZC9HXN29L9Ouoo8dZ3aS2HCYWQWLpk3TzL9p
GndtlwE1nWVv32wDNPTqbPTXJ/z8iVcRenXf9V+W7n7oj3vovlFkSqY5LprALd7I
8qrepAlEmWxT6HHc9LRPPRuxTCVBI0tSYa07ELUGKYW9GQUPK6xYhH5/AZUTzHVx
yKLKKhScNS1X56D3qjxQT5dJCbSG7GZl/3986kt/ALX1QGA/3cn0xt6tVtw3Ln8V
e1JRy1EZYm2kLvw93eAePT91u7RuRzeD9kU7GFoIFocscvo05vWqROyYA6tK8B4d
mWPlziSayQoDxMZS5ceaWZip5mweFaLM3s8PyNYPZYD11o/XnqNwWQqgNIf3UmHu
ZsaEXpCs+KpaBFt8WPmPXuymBfTTW6WxV67tNoAKRvLq1HS1i2CfAMrXhLZcuceC
d/WJjJWKyhofcvJbWWP42OdUWZd8pOJtRnzvdf2aBoUynH2pIub3kXJ4M13uX8jf
p75ApT0FUW6HW0tdzy3+GgBJey9vlwV0MlMCUfpDGK3zXNWSB0PBeXxRPW8MRjtl
kUS2SVsGVHpTNqxHtlHFl3rT8k+SvFxhkqQhkHByeB6so4P0asTJOad9vDZuyvxO
ViFdbRYiTVaN9Kf6JeYXF7VDIz0fW/PKaMnA0w+ZGihxvRxfmArLmejOIpvO8S3I
jjkp2HA4EU8YH7ovRVnUfLTABr0RZzFw/1sT3diHhJ5wvMkMQeTIoEvWxect3qMC
cZvofkNawyThcLKpJXv2FkAvKBRtEy2I8qg0yQnVSscA8l53Evdn2SshR2ZlTMDn
1CCkt6Pq5kgaKhXkeBR+u0MZWxnOQ7rjYYVL9i921LqUqb7/P8ipP6xw2S4e7Gfb
laC86F/Aoz2veU8QNZO9O5NQ1tRHYbzL+I7a46Jo7ORmD+yOkYOdDn/l+Kn6nYlm
4UXkLLVaRVX4ebpx97rR9GMnnOeQkiGcvn1RCFgSR06g+Gefcz+vldGNAcrAK2bw
5XjQLytXAAbMPZZr8TOH60vXLDlK+E+QKeabVngyWcHy6/91bgK5FJ09DJsQjwmq
fK704Dd/9CkjDKDZF3n8CNVZXuSkTJ6ZjjMtAl0aLZ0aq+ionyhim/fYJYbWtZ25
6oSZEMPes1tv736m6QQmkNCsuegdFvM3brreVaiX2MLZxC8snWaPwD7AYZg/45BZ
Gq077p49RWUsvLmgM1lSvAC7dpNbYQ+kdXUcR02IQx36bgR9Fk5pV5RThHoso4Y+
4XzLZB3pVWgbRFGTU3ThLvfq3bL/zH8LC+O1Jmb++71gbIcdyXJq5cdRSKLDs2g8
aWlqWrNcHCrWjTXn8wN59+ob4KGeIbWBvum8+eBg+AR0lfrFUOPIDfl/zQ+IRD2+
6agVQhmLX2KqcqxCy4LrP6N0XlhgcWUOSV33bXLspdZ9GCdQxHlnQE/2W9NYgm7e
jDqcl+h6tEuSA9yBc7cSBDGjuNLc/XbGTBGmN0V4iVGwKKyWWLmQn4cuMGReeYPq
hhQwUUrHUUPNBvqUprD9HLN4J0k/UH172N9tCo1jixddbWf39LHj1dvqAIsCXaU+
yv5Mpy0VHyWbIdutW1N/gfda7Dxk4aeurNTLwR16Ph21o61F69x44D11GSy+XDcY
oHxnmgK0dWjEPPH5oGXYU6QPC51TKoFbJZuIGZxlEBI9CZJfeDxCt36G+fOaDvaE
V5zw8Sl6CA50epbI9Qw609yivoGzX680oD7IXtpCn6KEhmEMWwCgBame5AIMeWVZ
kfSudn229z/mF0PKB8ELMNE1TyB5oQ2NUMTYfV7cEURVl5nFDRdRTk/tSp3EjMNc
o7NfeDhiCfMm8AFJSHpQRCUItJQShvNru38JRYAtYArT/IJ+MClAcPax3g8gmqmd
JnXc61Azo6J5JaepX5gCmJ7tVFqvcx4WhmuA33Lj3fkwhYGFUzLB+CZfxEMqmvg/
Qt/clg7InDK/WtnJbjy2DAsMGC98TFfzWteS/fHpvMmgvTHbOnWw3lFiVo6WdwZT
3bMYyCSsBWYtbZrVsFCD5sP1dK5Ip/49ftmJy6u2OXW8hxZD3MnyLxqVeIwRfbjo
QSgK3bMsUJckuBM6Xiw0JCghfXcT1drYHpwo7OlGmNAu+H+qea4Eex6rt6MXfGB2
ZyfZ3JhWJQQLXzUvNSH5DfyvIphAItboQC/U/GCb3fs/lIUw5oF3gh7At8fH7Kjf
0HJbXaY8tO4I5mggyF3KCNYqtMzBVNBWcFaxOjkrrVj7j0TnUMMxzHXqlUuvtbnB
cNXVHTzYqPWhyT4oICzidOLCorG1AFpGzcU/BPGrmWAEHEmmeg4PboecXee3J+jh
lDpt5QWmOCXizUYiZNRzQ6C6w3NVy14YrRoEpngrmmDsWkz412c3CAwUU6sp+tBH
s40iWdhgOBXAwiHEd6Tp7G1veNwyRFnRSTOWKpVZhW+ix2oSVqRaXInUuQL21PTr
sp2RKmpqcX0nFEJ4LyQEgZKGqp5Vxfy5D69PvfyQv6EUz1cwwLW/+YEy1CdQcf9q
DiAoMchWM9vgREZELHDz7PE4w4y0S+1DoN4gGB9ih1BIWZ2SixQRdreUKEviPA1C
sKDdE8+GtEn9ve8/xFJOun762/PiZ0UN0o8jwf94pUtrKGOM4hCwetd4uqid9Rma
WuksDecu2pXj/4iELjzP8gLCqaufLbtLteY/pac+PZk1yLUTDGy+NVn82N5Caugd
fMHEyyoeDtGIm8IipCtWLy9lidIY44+iDyclk++JWgYi08+dZoXpchB7OKSh4RFy
0I1sBwN55pCn8pPWvuDwjGL2cLx/9V4ugJ0ca0T8ekzD3MXvwLaQJPtyDJLQ2Shi
k/l2QlFRSqq9VkTU0zBiflHZt98nvH2eKwlfQJW2BDWYyD6giD6I+vVIzq9daTB8
694w43p6qL5oXZnVZ7RG1a1SWnKTtL5J7J+qSg1mPJAczC/S8DMHTEMiri2ryCg0
Q7Z2i+uFVMbIuQpqP+TAkElG/xxSWASM5buYJfn+jsedgaKDd2i4iNlToG0bOhCK
m49soPSqHNyv0BF9DchD7V0M1e5vTXRBbRvXEmN8c0BIXF5lvtFPeCliTtt7azNw
KpQ+NDlcxsL4OJBoehzZ7W7Sls8m8aReyPlDQxUE1WWrurYL0qXiMWL45on5N6XW
VkhE1cidIGz3QkqxT+PvxaIfZ1RgEWPhgl6wlIImYL8zFWaEva6JVSdL23Gcm0bg
HuIxEXeYhunP9HJeh0wry/PO0eL9ndQFDJynSvlQGUUbyYpee9bekAS7tQQA2tiV
JZIomY4OV3JySxk53VtBvF6ItpPVYtmZOnDw7B4RmuFOcN4N6qGZXJxWk+/iQ69K
jZkR4CZ31njGwlzuB7B9UG1dJuUVpSfLsMbkAekmy+MUouAIquZTlyWFzGVeaX5J
h0ec1Zj5mmnZi61n2IkEW0e8uICqHWv75EHxIzvs8KYnArhdTtgeyMZMVZnH5PIw
WVDRe8qDkNiUSXw5NQoSfPA0h+cAUa1bGhQh/BsB+0z2Mm4KewZw8sBAyrLObK+V
N6LQxiVzwcZ8pvuZN6sdBB0bz3uJMQicPcI8CQNJLgFQ+V3NFFArrw27JYIgYbAF
Fh4JpnPZKeokLsRkp2sRGn9cucK74Z0foXIEFSk7ovYIMeU/o06NfGIBaK0kX2VZ
SKJFamfNfiiagc/dpj96sgmuyQBWH05lJ5XCZQScx76JU//p29qtqCqcPL6LmKdD
DCtKWQNswKGiWYjIG9THbvGVVvs9WprzNFcedwCWqQORaxYaxtFv6n8igm83kfa9
0Zcb4I4XHIud+i8hCM5Snl1ruVBWxl0bswtI19QKb8U4fTyhpPMGdkseCbQ809lN
+lzWkPsrKQj0JN/iNzrMPegMKSXJjVGulr4sHjkyjz3NfZbGgyu66jDd0MsBvOU6
G/diEhEBDrTrGLO5/B08xLb/82vNZRxfF5MyL9A8HoGJk+ouGh0tzkYbY3tE1Xtl
kBTUMkwM9kskpwNLU9ugubf/oIBbKJyT5bogGv332vl5MnHar3ssYzz1WOcsX3lQ
ntBe3FuLQnjwlZTCOU9CowU4SHZDPFJIq8z+9VukvRBF01XAJ0P/h+xbKOFkbEBu
gR28yTbKzdP8/gAYaR1Z3zCk+HQHcUflaE+AtyGnh2hXWKhsGP1yB5LxaRrCfEsV
SbNzDtb77WS1CQYLpoVIYFxhL3HfUPdQOpfcs7x4YXZEOEHGRttuo8TBcLhtPDjT
hA7EsErYqJLw0eZFncMfFeX3yBLck5WPCHPGaSHrs1QrOYh6TfSKwvxvRfDEXinF
CA8olyyM4DOUve/9URdUa5571Ow7uzC433LCC3uPEGrxHFJGIMvCfRTPCCv7Cy8j
UwSC/lMdvc6f2M3xjerBtidUznWcjsMu+HZvrifK/IqmBvkIT7GQ7t+TbwX/ghqJ
zYBJYTwdd3QPbWXovTQ7bDD2/KcRyymQNZaSEC6Wiu6CwD4vA/peuMHoZVD/ShPL
xEOsEcGTJkelHdHSfqb32CmACHhU96re5orB3fxa21uxlMUZSHLoNR9YLmHacnLk
uWs8tPNJKYDZpRty2jpFp/I973CoJHRqpIUYxyTnX8wEwu0AamA8/cx+yQNk3Mfp
o6wIPTetmCyOT2ZSxWfD0ND6af/HOjNU6iVaU+dqaGQgHwBR0xpvBTUuHur7AL9B
LOCxdrIibfFtH/4cz3CeMGK+T3Wzp4eX/EzcAbFSo9FdSYNseof5hn/q1NW1Dyp7
FwnEabByz+cKm7y6v4cSsydROCCOcq2zHhAbv6uaRYY3dd5nQVE2WFPOy3rT3ayd
xmwHGiXjcU869cCHUehZwYysRBfj1miUlH91NVubDvXUAe/skBBgAdme0x2Njy4L
YcnbiTykvR4CrK1PnEa7eQ==
`pragma protect end_protected
