// megafunction wizard: %PARALLEL_ADD%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: parallel_add 

// ============================================================
// File Name: addeeer.v
// Megafunction Name(s):
// 			parallel_add
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 17.0.0 Build 595 04/25/2017 SJ Lite Edition
// ************************************************************

//Copyright (C) 2017  Intel Corporation. All rights reserved.
//Your use of Intel Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Intel Program License 
//Subscription Agreement, the Intel Quartus Prime License Agreement,
//the Intel MegaCore Function License Agreement, or other 
//applicable license agreement, including, without limitation, 
//that your use is for the sole purpose of programming logic 
//devices manufactured by Intel and sold by Intel or its 
//authorized distributors.  Please refer to the applicable 
//agreement for further details.

module addeeer (
	data0x,
	data100x,
	data101x,
	data102x,
	data103x,
	data104x,
	data105x,
	data106x,
	data107x,
	data108x,
	data109x,
	data10x,
	data110x,
	data111x,
	data112x,
	data113x,
	data114x,
	data115x,
	data116x,
	data117x,
	data118x,
	data119x,
	data11x,
	data120x,
	data121x,
	data122x,
	data123x,
	data124x,
	data125x,
	data126x,
	data127x,
	data12x,
	data13x,
	data14x,
	data15x,
	data16x,
	data17x,
	data18x,
	data19x,
	data1x,
	data20x,
	data21x,
	data22x,
	data23x,
	data24x,
	data25x,
	data26x,
	data27x,
	data28x,
	data29x,
	data2x,
	data30x,
	data31x,
	data32x,
	data33x,
	data34x,
	data35x,
	data36x,
	data37x,
	data38x,
	data39x,
	data3x,
	data40x,
	data41x,
	data42x,
	data43x,
	data44x,
	data45x,
	data46x,
	data47x,
	data48x,
	data49x,
	data4x,
	data50x,
	data51x,
	data52x,
	data53x,
	data54x,
	data55x,
	data56x,
	data57x,
	data58x,
	data59x,
	data5x,
	data60x,
	data61x,
	data62x,
	data63x,
	data64x,
	data65x,
	data66x,
	data67x,
	data68x,
	data69x,
	data6x,
	data70x,
	data71x,
	data72x,
	data73x,
	data74x,
	data75x,
	data76x,
	data77x,
	data78x,
	data79x,
	data7x,
	data80x,
	data81x,
	data82x,
	data83x,
	data84x,
	data85x,
	data86x,
	data87x,
	data88x,
	data89x,
	data8x,
	data90x,
	data91x,
	data92x,
	data93x,
	data94x,
	data95x,
	data96x,
	data97x,
	data98x,
	data99x,
	data9x,
	result);

	input	[127:0]  data0x;
	input	[127:0]  data100x;
	input	[127:0]  data101x;
	input	[127:0]  data102x;
	input	[127:0]  data103x;
	input	[127:0]  data104x;
	input	[127:0]  data105x;
	input	[127:0]  data106x;
	input	[127:0]  data107x;
	input	[127:0]  data108x;
	input	[127:0]  data109x;
	input	[127:0]  data10x;
	input	[127:0]  data110x;
	input	[127:0]  data111x;
	input	[127:0]  data112x;
	input	[127:0]  data113x;
	input	[127:0]  data114x;
	input	[127:0]  data115x;
	input	[127:0]  data116x;
	input	[127:0]  data117x;
	input	[127:0]  data118x;
	input	[127:0]  data119x;
	input	[127:0]  data11x;
	input	[127:0]  data120x;
	input	[127:0]  data121x;
	input	[127:0]  data122x;
	input	[127:0]  data123x;
	input	[127:0]  data124x;
	input	[127:0]  data125x;
	input	[127:0]  data126x;
	input	[127:0]  data127x;
	input	[127:0]  data12x;
	input	[127:0]  data13x;
	input	[127:0]  data14x;
	input	[127:0]  data15x;
	input	[127:0]  data16x;
	input	[127:0]  data17x;
	input	[127:0]  data18x;
	input	[127:0]  data19x;
	input	[127:0]  data1x;
	input	[127:0]  data20x;
	input	[127:0]  data21x;
	input	[127:0]  data22x;
	input	[127:0]  data23x;
	input	[127:0]  data24x;
	input	[127:0]  data25x;
	input	[127:0]  data26x;
	input	[127:0]  data27x;
	input	[127:0]  data28x;
	input	[127:0]  data29x;
	input	[127:0]  data2x;
	input	[127:0]  data30x;
	input	[127:0]  data31x;
	input	[127:0]  data32x;
	input	[127:0]  data33x;
	input	[127:0]  data34x;
	input	[127:0]  data35x;
	input	[127:0]  data36x;
	input	[127:0]  data37x;
	input	[127:0]  data38x;
	input	[127:0]  data39x;
	input	[127:0]  data3x;
	input	[127:0]  data40x;
	input	[127:0]  data41x;
	input	[127:0]  data42x;
	input	[127:0]  data43x;
	input	[127:0]  data44x;
	input	[127:0]  data45x;
	input	[127:0]  data46x;
	input	[127:0]  data47x;
	input	[127:0]  data48x;
	input	[127:0]  data49x;
	input	[127:0]  data4x;
	input	[127:0]  data50x;
	input	[127:0]  data51x;
	input	[127:0]  data52x;
	input	[127:0]  data53x;
	input	[127:0]  data54x;
	input	[127:0]  data55x;
	input	[127:0]  data56x;
	input	[127:0]  data57x;
	input	[127:0]  data58x;
	input	[127:0]  data59x;
	input	[127:0]  data5x;
	input	[127:0]  data60x;
	input	[127:0]  data61x;
	input	[127:0]  data62x;
	input	[127:0]  data63x;
	input	[127:0]  data64x;
	input	[127:0]  data65x;
	input	[127:0]  data66x;
	input	[127:0]  data67x;
	input	[127:0]  data68x;
	input	[127:0]  data69x;
	input	[127:0]  data6x;
	input	[127:0]  data70x;
	input	[127:0]  data71x;
	input	[127:0]  data72x;
	input	[127:0]  data73x;
	input	[127:0]  data74x;
	input	[127:0]  data75x;
	input	[127:0]  data76x;
	input	[127:0]  data77x;
	input	[127:0]  data78x;
	input	[127:0]  data79x;
	input	[127:0]  data7x;
	input	[127:0]  data80x;
	input	[127:0]  data81x;
	input	[127:0]  data82x;
	input	[127:0]  data83x;
	input	[127:0]  data84x;
	input	[127:0]  data85x;
	input	[127:0]  data86x;
	input	[127:0]  data87x;
	input	[127:0]  data88x;
	input	[127:0]  data89x;
	input	[127:0]  data8x;
	input	[127:0]  data90x;
	input	[127:0]  data91x;
	input	[127:0]  data92x;
	input	[127:0]  data93x;
	input	[127:0]  data94x;
	input	[127:0]  data95x;
	input	[127:0]  data96x;
	input	[127:0]  data97x;
	input	[127:0]  data98x;
	input	[127:0]  data99x;
	input	[127:0]  data9x;
	output	[134:0]  result;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "MAX 10"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: MSW_SUBTRACT STRING "NO"
// Retrieval info: CONSTANT: PIPELINE NUMERIC "0"
// Retrieval info: CONSTANT: REPRESENTATION STRING "UNSIGNED"
// Retrieval info: CONSTANT: RESULT_ALIGNMENT STRING "LSB"
// Retrieval info: CONSTANT: SHIFT NUMERIC "0"
// Retrieval info: CONSTANT: SIZE NUMERIC "128"
// Retrieval info: CONSTANT: WIDTH NUMERIC "128"
// Retrieval info: CONSTANT: WIDTHR NUMERIC "135"
// Retrieval info: USED_PORT: data0x 0 0 128 0 INPUT NODEFVAL "data0x[127..0]"
// Retrieval info: USED_PORT: data100x 0 0 128 0 INPUT NODEFVAL "data100x[127..0]"
// Retrieval info: USED_PORT: data101x 0 0 128 0 INPUT NODEFVAL "data101x[127..0]"
// Retrieval info: USED_PORT: data102x 0 0 128 0 INPUT NODEFVAL "data102x[127..0]"
// Retrieval info: USED_PORT: data103x 0 0 128 0 INPUT NODEFVAL "data103x[127..0]"
// Retrieval info: USED_PORT: data104x 0 0 128 0 INPUT NODEFVAL "data104x[127..0]"
// Retrieval info: USED_PORT: data105x 0 0 128 0 INPUT NODEFVAL "data105x[127..0]"
// Retrieval info: USED_PORT: data106x 0 0 128 0 INPUT NODEFVAL "data106x[127..0]"
// Retrieval info: USED_PORT: data107x 0 0 128 0 INPUT NODEFVAL "data107x[127..0]"
// Retrieval info: USED_PORT: data108x 0 0 128 0 INPUT NODEFVAL "data108x[127..0]"
// Retrieval info: USED_PORT: data109x 0 0 128 0 INPUT NODEFVAL "data109x[127..0]"
// Retrieval info: USED_PORT: data10x 0 0 128 0 INPUT NODEFVAL "data10x[127..0]"
// Retrieval info: USED_PORT: data110x 0 0 128 0 INPUT NODEFVAL "data110x[127..0]"
// Retrieval info: USED_PORT: data111x 0 0 128 0 INPUT NODEFVAL "data111x[127..0]"
// Retrieval info: USED_PORT: data112x 0 0 128 0 INPUT NODEFVAL "data112x[127..0]"
// Retrieval info: USED_PORT: data113x 0 0 128 0 INPUT NODEFVAL "data113x[127..0]"
// Retrieval info: USED_PORT: data114x 0 0 128 0 INPUT NODEFVAL "data114x[127..0]"
// Retrieval info: USED_PORT: data115x 0 0 128 0 INPUT NODEFVAL "data115x[127..0]"
// Retrieval info: USED_PORT: data116x 0 0 128 0 INPUT NODEFVAL "data116x[127..0]"
// Retrieval info: USED_PORT: data117x 0 0 128 0 INPUT NODEFVAL "data117x[127..0]"
// Retrieval info: USED_PORT: data118x 0 0 128 0 INPUT NODEFVAL "data118x[127..0]"
// Retrieval info: USED_PORT: data119x 0 0 128 0 INPUT NODEFVAL "data119x[127..0]"
// Retrieval info: USED_PORT: data11x 0 0 128 0 INPUT NODEFVAL "data11x[127..0]"
// Retrieval info: USED_PORT: data120x 0 0 128 0 INPUT NODEFVAL "data120x[127..0]"
// Retrieval info: USED_PORT: data121x 0 0 128 0 INPUT NODEFVAL "data121x[127..0]"
// Retrieval info: USED_PORT: data122x 0 0 128 0 INPUT NODEFVAL "data122x[127..0]"
// Retrieval info: USED_PORT: data123x 0 0 128 0 INPUT NODEFVAL "data123x[127..0]"
// Retrieval info: USED_PORT: data124x 0 0 128 0 INPUT NODEFVAL "data124x[127..0]"
// Retrieval info: USED_PORT: data125x 0 0 128 0 INPUT NODEFVAL "data125x[127..0]"
// Retrieval info: USED_PORT: data126x 0 0 128 0 INPUT NODEFVAL "data126x[127..0]"
// Retrieval info: USED_PORT: data127x 0 0 128 0 INPUT NODEFVAL "data127x[127..0]"
// Retrieval info: USED_PORT: data12x 0 0 128 0 INPUT NODEFVAL "data12x[127..0]"
// Retrieval info: USED_PORT: data13x 0 0 128 0 INPUT NODEFVAL "data13x[127..0]"
// Retrieval info: USED_PORT: data14x 0 0 128 0 INPUT NODEFVAL "data14x[127..0]"
// Retrieval info: USED_PORT: data15x 0 0 128 0 INPUT NODEFVAL "data15x[127..0]"
// Retrieval info: USED_PORT: data16x 0 0 128 0 INPUT NODEFVAL "data16x[127..0]"
// Retrieval info: USED_PORT: data17x 0 0 128 0 INPUT NODEFVAL "data17x[127..0]"
// Retrieval info: USED_PORT: data18x 0 0 128 0 INPUT NODEFVAL "data18x[127..0]"
// Retrieval info: USED_PORT: data19x 0 0 128 0 INPUT NODEFVAL "data19x[127..0]"
// Retrieval info: USED_PORT: data1x 0 0 128 0 INPUT NODEFVAL "data1x[127..0]"
// Retrieval info: USED_PORT: data20x 0 0 128 0 INPUT NODEFVAL "data20x[127..0]"
// Retrieval info: USED_PORT: data21x 0 0 128 0 INPUT NODEFVAL "data21x[127..0]"
// Retrieval info: USED_PORT: data22x 0 0 128 0 INPUT NODEFVAL "data22x[127..0]"
// Retrieval info: USED_PORT: data23x 0 0 128 0 INPUT NODEFVAL "data23x[127..0]"
// Retrieval info: USED_PORT: data24x 0 0 128 0 INPUT NODEFVAL "data24x[127..0]"
// Retrieval info: USED_PORT: data25x 0 0 128 0 INPUT NODEFVAL "data25x[127..0]"
// Retrieval info: USED_PORT: data26x 0 0 128 0 INPUT NODEFVAL "data26x[127..0]"
// Retrieval info: USED_PORT: data27x 0 0 128 0 INPUT NODEFVAL "data27x[127..0]"
// Retrieval info: USED_PORT: data28x 0 0 128 0 INPUT NODEFVAL "data28x[127..0]"
// Retrieval info: USED_PORT: data29x 0 0 128 0 INPUT NODEFVAL "data29x[127..0]"
// Retrieval info: USED_PORT: data2x 0 0 128 0 INPUT NODEFVAL "data2x[127..0]"
// Retrieval info: USED_PORT: data30x 0 0 128 0 INPUT NODEFVAL "data30x[127..0]"
// Retrieval info: USED_PORT: data31x 0 0 128 0 INPUT NODEFVAL "data31x[127..0]"
// Retrieval info: USED_PORT: data32x 0 0 128 0 INPUT NODEFVAL "data32x[127..0]"
// Retrieval info: USED_PORT: data33x 0 0 128 0 INPUT NODEFVAL "data33x[127..0]"
// Retrieval info: USED_PORT: data34x 0 0 128 0 INPUT NODEFVAL "data34x[127..0]"
// Retrieval info: USED_PORT: data35x 0 0 128 0 INPUT NODEFVAL "data35x[127..0]"
// Retrieval info: USED_PORT: data36x 0 0 128 0 INPUT NODEFVAL "data36x[127..0]"
// Retrieval info: USED_PORT: data37x 0 0 128 0 INPUT NODEFVAL "data37x[127..0]"
// Retrieval info: USED_PORT: data38x 0 0 128 0 INPUT NODEFVAL "data38x[127..0]"
// Retrieval info: USED_PORT: data39x 0 0 128 0 INPUT NODEFVAL "data39x[127..0]"
// Retrieval info: USED_PORT: data3x 0 0 128 0 INPUT NODEFVAL "data3x[127..0]"
// Retrieval info: USED_PORT: data40x 0 0 128 0 INPUT NODEFVAL "data40x[127..0]"
// Retrieval info: USED_PORT: data41x 0 0 128 0 INPUT NODEFVAL "data41x[127..0]"
// Retrieval info: USED_PORT: data42x 0 0 128 0 INPUT NODEFVAL "data42x[127..0]"
// Retrieval info: USED_PORT: data43x 0 0 128 0 INPUT NODEFVAL "data43x[127..0]"
// Retrieval info: USED_PORT: data44x 0 0 128 0 INPUT NODEFVAL "data44x[127..0]"
// Retrieval info: USED_PORT: data45x 0 0 128 0 INPUT NODEFVAL "data45x[127..0]"
// Retrieval info: USED_PORT: data46x 0 0 128 0 INPUT NODEFVAL "data46x[127..0]"
// Retrieval info: USED_PORT: data47x 0 0 128 0 INPUT NODEFVAL "data47x[127..0]"
// Retrieval info: USED_PORT: data48x 0 0 128 0 INPUT NODEFVAL "data48x[127..0]"
// Retrieval info: USED_PORT: data49x 0 0 128 0 INPUT NODEFVAL "data49x[127..0]"
// Retrieval info: USED_PORT: data4x 0 0 128 0 INPUT NODEFVAL "data4x[127..0]"
// Retrieval info: USED_PORT: data50x 0 0 128 0 INPUT NODEFVAL "data50x[127..0]"
// Retrieval info: USED_PORT: data51x 0 0 128 0 INPUT NODEFVAL "data51x[127..0]"
// Retrieval info: USED_PORT: data52x 0 0 128 0 INPUT NODEFVAL "data52x[127..0]"
// Retrieval info: USED_PORT: data53x 0 0 128 0 INPUT NODEFVAL "data53x[127..0]"
// Retrieval info: USED_PORT: data54x 0 0 128 0 INPUT NODEFVAL "data54x[127..0]"
// Retrieval info: USED_PORT: data55x 0 0 128 0 INPUT NODEFVAL "data55x[127..0]"
// Retrieval info: USED_PORT: data56x 0 0 128 0 INPUT NODEFVAL "data56x[127..0]"
// Retrieval info: USED_PORT: data57x 0 0 128 0 INPUT NODEFVAL "data57x[127..0]"
// Retrieval info: USED_PORT: data58x 0 0 128 0 INPUT NODEFVAL "data58x[127..0]"
// Retrieval info: USED_PORT: data59x 0 0 128 0 INPUT NODEFVAL "data59x[127..0]"
// Retrieval info: USED_PORT: data5x 0 0 128 0 INPUT NODEFVAL "data5x[127..0]"
// Retrieval info: USED_PORT: data60x 0 0 128 0 INPUT NODEFVAL "data60x[127..0]"
// Retrieval info: USED_PORT: data61x 0 0 128 0 INPUT NODEFVAL "data61x[127..0]"
// Retrieval info: USED_PORT: data62x 0 0 128 0 INPUT NODEFVAL "data62x[127..0]"
// Retrieval info: USED_PORT: data63x 0 0 128 0 INPUT NODEFVAL "data63x[127..0]"
// Retrieval info: USED_PORT: data64x 0 0 128 0 INPUT NODEFVAL "data64x[127..0]"
// Retrieval info: USED_PORT: data65x 0 0 128 0 INPUT NODEFVAL "data65x[127..0]"
// Retrieval info: USED_PORT: data66x 0 0 128 0 INPUT NODEFVAL "data66x[127..0]"
// Retrieval info: USED_PORT: data67x 0 0 128 0 INPUT NODEFVAL "data67x[127..0]"
// Retrieval info: USED_PORT: data68x 0 0 128 0 INPUT NODEFVAL "data68x[127..0]"
// Retrieval info: USED_PORT: data69x 0 0 128 0 INPUT NODEFVAL "data69x[127..0]"
// Retrieval info: USED_PORT: data6x 0 0 128 0 INPUT NODEFVAL "data6x[127..0]"
// Retrieval info: USED_PORT: data70x 0 0 128 0 INPUT NODEFVAL "data70x[127..0]"
// Retrieval info: USED_PORT: data71x 0 0 128 0 INPUT NODEFVAL "data71x[127..0]"
// Retrieval info: USED_PORT: data72x 0 0 128 0 INPUT NODEFVAL "data72x[127..0]"
// Retrieval info: USED_PORT: data73x 0 0 128 0 INPUT NODEFVAL "data73x[127..0]"
// Retrieval info: USED_PORT: data74x 0 0 128 0 INPUT NODEFVAL "data74x[127..0]"
// Retrieval info: USED_PORT: data75x 0 0 128 0 INPUT NODEFVAL "data75x[127..0]"
// Retrieval info: USED_PORT: data76x 0 0 128 0 INPUT NODEFVAL "data76x[127..0]"
// Retrieval info: USED_PORT: data77x 0 0 128 0 INPUT NODEFVAL "data77x[127..0]"
// Retrieval info: USED_PORT: data78x 0 0 128 0 INPUT NODEFVAL "data78x[127..0]"
// Retrieval info: USED_PORT: data79x 0 0 128 0 INPUT NODEFVAL "data79x[127..0]"
// Retrieval info: USED_PORT: data7x 0 0 128 0 INPUT NODEFVAL "data7x[127..0]"
// Retrieval info: USED_PORT: data80x 0 0 128 0 INPUT NODEFVAL "data80x[127..0]"
// Retrieval info: USED_PORT: data81x 0 0 128 0 INPUT NODEFVAL "data81x[127..0]"
// Retrieval info: USED_PORT: data82x 0 0 128 0 INPUT NODEFVAL "data82x[127..0]"
// Retrieval info: USED_PORT: data83x 0 0 128 0 INPUT NODEFVAL "data83x[127..0]"
// Retrieval info: USED_PORT: data84x 0 0 128 0 INPUT NODEFVAL "data84x[127..0]"
// Retrieval info: USED_PORT: data85x 0 0 128 0 INPUT NODEFVAL "data85x[127..0]"
// Retrieval info: USED_PORT: data86x 0 0 128 0 INPUT NODEFVAL "data86x[127..0]"
// Retrieval info: USED_PORT: data87x 0 0 128 0 INPUT NODEFVAL "data87x[127..0]"
// Retrieval info: USED_PORT: data88x 0 0 128 0 INPUT NODEFVAL "data88x[127..0]"
// Retrieval info: USED_PORT: data89x 0 0 128 0 INPUT NODEFVAL "data89x[127..0]"
// Retrieval info: USED_PORT: data8x 0 0 128 0 INPUT NODEFVAL "data8x[127..0]"
// Retrieval info: USED_PORT: data90x 0 0 128 0 INPUT NODEFVAL "data90x[127..0]"
// Retrieval info: USED_PORT: data91x 0 0 128 0 INPUT NODEFVAL "data91x[127..0]"
// Retrieval info: USED_PORT: data92x 0 0 128 0 INPUT NODEFVAL "data92x[127..0]"
// Retrieval info: USED_PORT: data93x 0 0 128 0 INPUT NODEFVAL "data93x[127..0]"
// Retrieval info: USED_PORT: data94x 0 0 128 0 INPUT NODEFVAL "data94x[127..0]"
// Retrieval info: USED_PORT: data95x 0 0 128 0 INPUT NODEFVAL "data95x[127..0]"
// Retrieval info: USED_PORT: data96x 0 0 128 0 INPUT NODEFVAL "data96x[127..0]"
// Retrieval info: USED_PORT: data97x 0 0 128 0 INPUT NODEFVAL "data97x[127..0]"
// Retrieval info: USED_PORT: data98x 0 0 128 0 INPUT NODEFVAL "data98x[127..0]"
// Retrieval info: USED_PORT: data99x 0 0 128 0 INPUT NODEFVAL "data99x[127..0]"
// Retrieval info: USED_PORT: data9x 0 0 128 0 INPUT NODEFVAL "data9x[127..0]"
// Retrieval info: USED_PORT: result 0 0 135 0 OUTPUT NODEFVAL "result[134..0]"
// Retrieval info: CONNECT: @data 0 0 128 0 data0x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 12800 data100x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 12928 data101x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 13056 data102x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 13184 data103x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 13312 data104x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 13440 data105x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 13568 data106x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 13696 data107x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 13824 data108x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 13952 data109x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 1280 data10x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 14080 data110x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 14208 data111x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 14336 data112x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 14464 data113x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 14592 data114x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 14720 data115x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 14848 data116x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 14976 data117x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 15104 data118x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 15232 data119x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 1408 data11x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 15360 data120x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 15488 data121x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 15616 data122x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 15744 data123x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 15872 data124x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 16000 data125x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 16128 data126x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 16256 data127x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 1536 data12x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 1664 data13x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 1792 data14x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 1920 data15x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 2048 data16x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 2176 data17x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 2304 data18x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 2432 data19x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 128 data1x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 2560 data20x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 2688 data21x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 2816 data22x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 2944 data23x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 3072 data24x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 3200 data25x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 3328 data26x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 3456 data27x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 3584 data28x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 3712 data29x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 256 data2x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 3840 data30x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 3968 data31x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 4096 data32x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 4224 data33x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 4352 data34x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 4480 data35x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 4608 data36x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 4736 data37x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 4864 data38x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 4992 data39x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 384 data3x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 5120 data40x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 5248 data41x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 5376 data42x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 5504 data43x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 5632 data44x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 5760 data45x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 5888 data46x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 6016 data47x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 6144 data48x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 6272 data49x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 512 data4x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 6400 data50x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 6528 data51x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 6656 data52x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 6784 data53x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 6912 data54x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 7040 data55x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 7168 data56x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 7296 data57x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 7424 data58x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 7552 data59x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 640 data5x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 7680 data60x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 7808 data61x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 7936 data62x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 8064 data63x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 8192 data64x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 8320 data65x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 8448 data66x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 8576 data67x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 8704 data68x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 8832 data69x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 768 data6x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 8960 data70x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 9088 data71x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 9216 data72x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 9344 data73x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 9472 data74x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 9600 data75x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 9728 data76x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 9856 data77x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 9984 data78x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 10112 data79x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 896 data7x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 10240 data80x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 10368 data81x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 10496 data82x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 10624 data83x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 10752 data84x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 10880 data85x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 11008 data86x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 11136 data87x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 11264 data88x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 11392 data89x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 1024 data8x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 11520 data90x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 11648 data91x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 11776 data92x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 11904 data93x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 12032 data94x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 12160 data95x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 12288 data96x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 12416 data97x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 12544 data98x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 12672 data99x 0 0 128 0
// Retrieval info: CONNECT: @data 0 0 128 1152 data9x 0 0 128 0
// Retrieval info: CONNECT: result 0 0 135 0 @result 0 0 135 0
// Retrieval info: GEN_FILE: TYPE_NORMAL addeeer.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL addeeer.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL addeeer.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL addeeer.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL addeeer_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL addeeer_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf
