// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 17.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
T+8dyVjZD4FtxuhfB9MLMobDws5vXx/5lgZK4QmpueKyy894bSFwd77Z1XuAetX35vcsBQxn6D2P
IxwmYsEcUVq++W3f3vX45L9MWgwRp0kNDHOxnmiocjJHyqhIVFWb+zPWDds8n4WFipHmKtdMLVjX
8oPbRZ0rYHMElSFpIqD0tRgTtKpR2+v2J0hu9KrJ0aqxlnVKc1SekiqydFzwAsQ4XfR2bQCYGQRJ
8qKcdF80iHFMIM6M0YjFvZ+sKEYKtpqBSw5PZMzuPM9kQceR5Ms6dwLvUGE/1iO3DiJJZXVooEAc
JHE3+1dIIsYsftJlxMMIhEUoqIgBW0LYfDdr0g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5760)
EylRTQquTDa+46xOML//OfI0JffNP7QqGqABbcRyNKVDEHmaj5kBI66u6hcjzTDlXXYAebkPJLud
avVQJ05hxG5OgdjvtH+UQ+ft01AXGBneTpCsrW9KfLg1VVFJvvNlyQDo4AXbXYvFWQP21Xud/oRv
q8j7u2gDeUbtMl6/O2vLTgOTTtaQ3X/aNy7199QN+gQxoWchxTBk34+cknCB5GhLP7ZsQ1PRAhBZ
1JiArHr1BhRD3hqLk6WOUeE2xAc3kioaEohRPlB1sUHg8ISCEvg0AUHixXBz1XWm3zIZA+Y2iPcN
08dpx3WIPGEHgHhq/TZMR+Stdk4NuRS3WPQHfykkmGCKWD7lG3X03sekq4CHJm8NXE/cc6S+cm1T
zjNb12u0gj/TSrVNrFkWVFv9H5tnqeXXCJifwBXKWANa7g59sA1mBczlzBSjj6lBVHk3DZWGQYVZ
fdim/HmJIOdFgJkGDS9pzrvoAGlVwtTwIBGTC2JzGUKUNdpwREfu2gT8azcqppC4iQT996SOAC97
2c+zQu9UfuoLw1p9IvBFNgDASXzr0Fe1/8FCV2OTPWdSNvahQkolznm6FCFrnWnpZIkLg3X7Cvx8
XpU8+IhsampxGoi1fJy5nl8gYcW8TMTUJEZKltRjSSBRGKrVkWcfQqynP0AGbLaqstYYn4XGUy7z
QjDs9oYZl7Ngd9EVcmwaDoPccgheav+iZqkocd90dg10vIpg1Ldk3EwN9stB5q8PXGpt9a8x+uX9
XRRUcwzDckMTpAKwKSwdPECZKPHpHVeS2bbbYdjSSN8dewYNJgj1pRu6CLfvQFObxDOM8JTyOFae
5DxrUEDtyCrZZzAGIsG1Y+YtbniEQzcBgfyJC/pTLxL7j3TjTodDFUdKbvTKSrhXvCIbsn7hMPLc
V8yAZkBrwHUK90FOh9uDxN2ibNl57GL3/lTxVirOnbwZcCcmL4r4af+rlm8AsLVT+7Yv3+SUyD9c
KnpGaNCL1x/bZ3cG+6NLYxyguUphvO4gqCIcigJR8Ql/3AMHRsmJ+XvbtaB2szSBMI0rT+xbizMz
bcmtK3c57/z35gjxtPlamdPMh3Yp2qYIcAJ8fUUsg/DvNidIVK9F60pdZDG3ls+ooTAOPIxODD9s
RpHbDt0/Ugc7+8q/NCHhXfcjoQInrwbPz+UH+3WSlsb98ruleE38htt+PG7xHTzFKgU4LGjbTMyV
0IqGeBNj9Co8xzw1eQPSQtzNnOzOLqJFam0YLrelULdLr3sGyd2IrQoOBOvuYuzuHvsiyr9RLto6
QM3xYMxmGcrZOOmat1LQpzFKF3jr7JnyxZWMETeGu22arlGcl+ucTeYxR7stSqYrZ9bzzcN5vWGD
2lmNbi/SePa1lM4kQcgwJMYH2g1Jv571e81fODZ09gThInFVQV5iXPPk2rsQqYSOX4B+Uite0YBM
A9JmRJchLt6yKaYqgZgUpwnKmSA1kRGNWCO3WSfAjFE3pVdVpgiughGvHw9XYE5m/ui1QZqLlEPt
+Ek+6EJ2gMHm9L3tIsqWh1ayLfdGbG2f3nlm1HauHMboJfh5x4FzkFvYrslM7iQE64JidER8dqmr
sJBQwWApBqZeO8bn7BzRqtgfRYdgTaXywIoJDJg69P5uRux4zdplplj5u3jwJBFGAAAoRYHTfg4Q
Ti+KnpYh+/GngCGa2RmAga0hPtVDZZhsoc5FZUI2Vdz+Q/IZ6tW5dl4W0GsITAG9RTk2koUM/Dd2
esJBd0ZGuwk3hq2zQqPXVYN3mKttjs1hikMGxjXJiywteWE+jRSzOfhMxeFM0R5OBnae/I0wC/36
SpVsUdbhbQfUll8w162krCK6TaBSszOhVjyAfet16zUFlFQoUaSq6abmrTm5cL9ksznLXcwk/iXb
Py9+cKjJUtl4GoxiwLCXjXCOv/NhdO0v2PnK3au0psbEW7v/NW5KdAEuiNIvAc+G6zDf9BRCpOzv
CvZwxHPXWVwUE340bRtVHKRJyI5EldGO6sjryIFs0+ZJuxCTFvqPb9vHZddCAbiaL5j8/qO2IhF3
fWHx69NRyAPXlg07zYZbU3P7hMRN6EGFORYv0spJC+9VRCuR1rwKlP2ONOyGWfaGZVZIEpyqsdgm
sYNlmsEEnnRrw6xNK7wGoZK8EePjOPniXo0fJawA8ZJ5zFerCUfuaV937CsjiOPc6JU4ERuBEe9r
Eftp1JSkvooovph4HZKyyzv57Ogwq3gisSABk6q2sDbdLXp3im1hX4esqbheElHfBQQlNFutdp4F
sC8FNRd8FN0dsJg+dYyqK9L8YxGw70kpGy8YJcjmYtBghKotBfAUzLClqnKZRJ1OXp1P/wFU0ZvW
ozANrmPrTeUDm/+kHTVan8EqZTBiuTO3fwEPF3wqvkNAnlqTT3+gxHOULiGZQYbpBxm8hTc7+CaK
QS7nHivDeNylbkQZKLDQbxFMS/LVqTqGxK4eFRLX84HIBm8olL1eFhE7zEHPlSEYs6Y2m63G1Vb4
eGyAVbNlhVJ0hOjvtSImLu977xLOdHk/BWFJSy15doAfyaOQv81Y0PuIusELBVW4M8om7GH7ZVD+
bpH8K0hnSaY62hN3MwcmegLLVose5FyICM1m1AE0U1vSXL/v5vou6XVLHaBjPujjcFLwuzRA2XiB
VYrDtqzJN2puDqfUi8efce+KsmRFKHz7ve4sLP75nlOkUZ5LJloA0WybRQV3gbuIo69VG9edvFrb
nWkxMw6WP70Ln61dGEwO9Tc5L/ITk0U1biOSIoMVgK+R3TL63PFkNYDosirC8wJH/ZqyEYyS4hZD
NxGMjeU8YI8zdzkTmJdecXD2bCxrTQAQBPqPoKTXwQZfIreKI0ewTSz1D+v+Q110b/M8NUNhJvr2
OgqqvpHkAYkn1AyS9e7ti2Gfl5SIsYmXOfifVGBikcAZXMrq6heztO/Qe9QRKcZVXTbloKlsiTk/
a/5F+63SdYb2mUyfipe40pr6TmGgvRm/EUvlTTOZOg8a+vH8uvD9uJcOt3ZymmJbj9aqBFxG6Kpo
7/EAu7EUQ1JRlL2e1E5rdfc9UBVlkm0c1W1IDidRvIQ6X0b3yiVpQWCXCeuh/VqnBj4xY0jrDM+D
EYj/83wmCnvPcYQtGNwx/K3llP7hZQpqFN6a3PER6Yf/cuYXtnDmTlREwx46Izuwzkd7H4NScTNW
XXMHjHEiSljl9yYiTtA+hAzWkNkRqzUNVKp19OPjXMPU4L9jeGVhW6rR4MzV7YkCZ+MpdZ2D8QxI
P5TmJAFkDGNd3Ne/9/FkTEGkscqUD6mJn+6lhafxY+FCmMdtMsUZnFnmxycIOh1BAT1NbLpNsQMf
r/6GWY7PG+la3/b1e9LAmGddlR0sNL14bFyxZEZIAyVWfWgTKZTAXsUzTkwIImS07NCD7p3ISie4
0hT1epTItAvLjCh7V+seTZXqZyjzdgGad80N6y7jNfKJfU+hwhu+NT4znMuBWXnn9ojKWsjdWuno
tuVruM6UU4WE+MY1D/cT6GV5OFBpaA+A165reUhgV/o+78osSb0RyO4CtnViKpmp2R3auZZgspGs
3H0Lyj0NeDFixN48/h1Ol4fyrGrJAKajL/YvyqaMjMlW8b5TMqdinXtWEJ7AJTLiXRyMFBm8ZUiW
G6TYoXRBjZLM7CnTuz92g2mvSzsdfN4pfpviT6KzH75tWpcr3TM3itd7ZLc+d9md5y2YfB7v5CWp
Vmr/0T8GtjaaAU4+arIb9q+j7OAVRdmO4tugCkKe8hxdhIk0BzD5Wn1rUO64CehVb9vRvxrY6DpC
/1xBz0+HtXoMrWZZ2cvj5lpPcsFxuOW5vqixXmeTzIqJCn38/SwJO96aQv0oU5HcZMTTD07+AIZE
JMb1tVfELgmh6/cn5hzYHOo3mvgrBV49L+ZOtlUh0GqqnnIyNbS9jVxXvulJyzIu5e6jcMRydAmK
RDFkIigLMDWjwkb2hrgeAsk5AuYYFPccJ2QX4IzLSm3DgNMwkB5UCzQnXrwxCnXkr00G9/x0viOR
8Mjo7/p8ANQGUGJ+TjdSHmchhwZ7kFPSyUmm5JigV/fiTfH51MzsbBIC8xWRbzrmO761Af8wOIH5
YC2vAMGwACP8X+Q+VidAkS/goy23kovUoWSQOm0s48k6PbzG6x0WlmobMWr+gB0wS3gUfYYwLDXk
vPID8MQuKjMKyTcjS+tfohN2rTtGZ6LZJUicYBZ4x6w05pU7ZdhOOAXs3pE2MAI5MEGggOOVoCdW
PcqA5Wnvy0OskgZdoQ81yYRvHQEO+jbiWrOI0W5NF4UEVBF3uG9Sim4AkcocY8X7cmxvQ8r9nlBc
EpmdO11GAoYI2jRHxOwTNqaAwJiM5GVSmLi5rvuVrrAzxGXMtaqMluyrrthOzqdpeNpuCo2oocsf
YM0rDYj7Gq2Ix3Jjh1c2yvLtf4bxItsv6uFJAtz2j7ji+46GKFe9WHxw4aHVkgY1Vy1K+p5YtT6O
ztMbONDVEM5qEPgH9bWm1iwNGLwq0t5FnMuQP0gthIf6siTnWZ5NHtEPArrZcZiiSTcPhqoUD1QW
Var54e/FpPY+ovXENpBK6zwKZV+KY96Z8KcdWAdR/yv5ywlG5X1ug6MFwr7fc3Fiv33GgSn4wLsZ
rAz8Xyo24jNeZYrYN1w8t5SWxJSzFDwmO7MqfCjZhKg/fObwasmhYWLB8tsD4o+ppfFqviKHH/vW
MA0nVo7V1qKFyPmhimQDRolJFHyY7VQhHGeWcKdw+F7WX37M22WSOC3FFc2ItODop5HcVBh9x5vc
NhKpVvaZPdzSbrkmlGZyek/vbSi6BD8EqveMs+fpp7HWrRCEZ8ey2bKk9jHnynZ3fT25MRVPIaGc
AVPgJCTVnY6LMUExuq0KQmTPJ0D4ba7UzCNoTeXNkWeT++X0+N8MfMFMCBdBRlBAszgls8NXTV/Q
AlGj4eMt0m8XH4fWfFX1m7WnCW905H7j6l4Rs8dxd5Ij2iUloFHn27k2rd1amEWDKl52ubfjj9zc
kKynGM3mfVOszxBZ7pc+Z7bLkXM1hl2HOmy3pjR2D7g3bPXqhEBx+g2M9YfAWY9QV0yGbBqHmbNn
CR7OfsVTLozqCnaVa9g1Os90AWVluZZ0jWWH3oKodDPAsi5FU9VNM1cMUh9AElW/sDB4jKTxRPQw
0d6CuJKHd73PhUFnhsOOiz5JEy4XPZZ3Hp6MWSnlITnbV4JqccMnIQ4IC/o3hdNo6kCsI0agZ+MC
jGkhD4nz7R2Qg48fTdaji29UDbLoDOOjYQQF7SxlCqrd8FfvIk4Z4Rb1EXliDB98+oGZ8bVqcf4x
QzpOBtQuXil488b3a68nVdCbziCqDwP0a6w3HrRWTpbz3ga3DKti5zSrWKZmN5A2sOdDCqBlgTXt
7uz/UzP7GfnzC2XhweAHkgdFgbCO7F0kzuJ2FSBUjkVR5fN23+qOzzJ31gRWbPFz/Mj18fQBrY+w
x4Eu1BpeJDGCGl9MmLqnLeyBVydN6rpXHn7H/zmEcBHgLhyqrPQCbXaJhfSySnPWVQQliyt4ok1e
tCetcApJiGvtmajial0VLuoGmHnyAS2jGzErYIAz2eNAb6NkfHXHhbnQncKKpOebOwUlPn0NyMrz
B4ZuN1iLf7K4POzkPtOPajInjs2jnErjYYMjYlMq0CJbfiBDuN2soOH1n8ESQMt9rTqvLuO3DGnL
qNhkcqNsGfyHaorfoRI72qw21HN6RNYYwUUHcJnJq3WOHODXThSxUcb7g7PzbTccKSdlmpaSsR8f
LzhruhURyr3JCtzBORKsrHyx8rj9hLJQvoc4oU1H1tJQhrRcHyBR/GPrODruf/jO5xG7nWCZBJNs
olfraqh5ict4i37BKFbN+uoCLH0E8I+ZIwg2ygVzLRwlB2FsLGzhb93s1PQeS9psuxVLaPegPO3/
DbTaYLVOLakSZGJX0KBrCgGhhHRTYyvEdTOON+dUw6jLki8fjWmZa4hgbthrYaY3EyhkSQ93d2+6
C9qfvQeY4xqJhreyNM+wsmum6Op6EgzjVhLkq/bZ1s+hgE/54hCgrJRBVdvyS9mkGaqFb7PIhmW0
qcrOBXmoMqMTXJJeofjw3urVQkRMazQm5IKVK62yLZjywqOPw5jomI8XqAsH1tATzUkSUTf+U0qO
gVBGfs03vo6lgtLKtiWguUl47d40dSAaKVMDdmalTBupwjyBwY7MBmGUqTCiVuZ07pcc5vlMj5Z3
OTDOWA+Ivqn3y/5vdmZO3bJMc4ihi7DZqqX52CszpZrzhsbacBN9EAtZgKhYlMm+i9MP6T7RBTko
AdnIJusApWJag8oTeJXCcPmkGdhJh+D1M0IiEN8VVBnVeD9Orp8PUQkY+29SmKTDg9ZlRquSmDbo
z3pFtD87pmSjavwTImpWXFpNDOTUIwsGiBEOCV4E/6KUsgmrJ4i2QGwvfOQKmDUdbc8QQXQHzwlt
67mmVeIV7JtrD9vOnVEUcyE9gFbXVIk4owEwmpER6y/uT83QRVpXNWKFluAERndf4JrpSMqbxEEk
6Z2rdsaZDiaxzRaLi26/NiyWxQ0M8W7+eO11nmCdYzlXNFbRcxuxQ684fsyudLecXqDceOBT92XW
Z4GZeWse5lvq0S0aokufuJ9MyqPxjLYcA21LZWKP1/WnB9ZsZovCw3nwTXMfLv292KI9x5QbJbob
yhjtmNYiin/Y4BzixEZC+ULedXTwroC55RZ3aJObSq5rcmnwcmSFjCTd+fqurvpsg4TT8/It/UHE
ilLGj7hKhwBbYI4AgFZavLxgou5iJoGd+eL9wUAUajC348ceNVcWfrzAKmVdnWGQA6TmlJBfrH77
Rqgjf1DKqfezkQkoWEbhPDuEjgaQ5gsawgf+zhvbhJhJBO3ssbTcoDLslozbTJX7FUm5eOzh05Qr
y2vYs1wz+nBrZXac9+FAONB+8zjYZkJLRPO/HT9eDvPIIBR8dzMHezebzJ6J5g4DdDL3wm+uLaWE
OGsfFEzZl3L0fVCfCG3Z1HtZTy68fRQmXbufrvAdPKINdGZnSim3IBg3IZGSdzTxdAwblcxJaPL2
KEyDY3ix6Lp2z+6i0zflZq8WEFCsmjJFcggzkV+Xq4rcyx3vn32g890NPN2WSosnvR+9yCt7XtTh
/moQ9zeKrModj4vhjy6ZHICciKH6amX3bqxWkriVK1Lz/onJ0KW0Go42VyyKetumeZwtPiTJu7u/
e7UstzYG91ctyL+eJFfCffgjimocyzJ2azlRUx2puB0DAlXaAMJvCaO8sOq0XeIsJkOe9VWiIoe8
8y9Xya90JQzhnUhqWKrnSy2vVDAHuyfldi6DHlP++nDzSuz56SGpVR6+afYPjLCVpSvypwAGoiNL
fAeDKeChIt0Uj8HmVD7ZGSd4B6yy/5S3hXp/qQWZR/ZKhtCNK5E2KlbIS+rdDNj3pIt59EP2Ejxa
SfrU365VqdXp581/U+VhUC7Fo81juHcuxXTf/h9tG7fRGKCe7RS5Cfjk7H8np2CKgSlQKq9jq86y
8+M6qTLdwaQUvTcFvxne3B1Gmh8hy7c5/LM7BGDZ3ajIJbsnPxYccK8u3OT1tsEglH85aZ2j/kYj
kM+B8OHQUSEFGniTp5Mbt2lnmKCtknRGHAqL40psvkPW63ExPsKhKbdmOO42ilaJPeO0PL1fPSS1
fz6c
`pragma protect end_protected
